module BOOT_CTRL(
    input   wire    [3:0]  state,
    input   wire    [0:0]  end_m0,
    input   wire    [0:0]  end_m1,
    input   wire    [0:0]  nWAIT,
    output  wire    [0:0]  latch_d,
    output  wire    [0:0]  rst_mb_addr,
    output  wire    [0:0]  inc_mb_addr,
    output  wire    [0:0]  rst_m0_addr,
    output  wire    [0:0]  inc_m0_addr,
    output  wire    [0:0]  rst_m1_addr,
    output  wire    [0:0]  inc_m1_addr,
    output  wire    [0:0]  CEN_MB,
    output  wire    [0:0]  CEN_M0,
    output  wire    [0:0]  CEN_M1,
    output  wire    [0:0]  nRST_CORE,
    output  wire    [0:0]  BOOT_END,
    output  wire    [3:0]  next_state
);

localparam ST_IDLE	= 4'd0;
localparam ST_REQ_MB	= 4'd1;
localparam ST_WAIT_MB	= 4'd2;
localparam ST_REQ_M0	= 4'd3;
localparam ST_WAIT_M0	= 4'd4;
localparam ST_REQ_M1	= 4'd5;
localparam ST_WAIT_M1	= 4'd6;
localparam ST_BOOTEND1	= 4'd7;
localparam ST_BOOTEND2	= 4'd8;
localparam ST_BOOTEND3	= 4'd9;
localparam ST_BOOTEND4	= 4'd10;

reg [15:0]  tmp1265807652120;
assign    {latch_d, rst_mb_addr, inc_mb_addr, rst_m0_addr, inc_m0_addr, rst_m1_addr, inc_m1_addr, CEN_MB, CEN_M0, CEN_M1, nRST_CORE, BOOT_END, next_state} =   tmp1265807652120;
always @*
    casex({state, end_m0, end_m1, nWAIT})
        {ST_IDLE,	1'bx,	1'bx,	1'bx}:tmp1265807652120  <=  {1'b1,	1'b1,	1'b0,	1'b1,	1'b0,	1'b1,	1'b0,	1'b1,	1'b1,	1'b1,	1'b0,	1'b0,	ST_REQ_MB};

        {ST_REQ_MB,	1'b0,	1'bx,	1'bx}:tmp1265807652120  <=  {1'b1,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b0,	1'b0,	ST_WAIT_MB};
        {ST_REQ_MB,	1'b1,	1'b0,	1'bx}:tmp1265807652120  <=  {1'b1,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b0,	1'b0,	ST_WAIT_MB};
        {ST_REQ_MB,	1'b1,	1'b1,	1'bx}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b0,	1'b0,	ST_BOOTEND1};

        {ST_WAIT_MB,	1'bx,	1'bx,	1'b0}:tmp1265807652120  <=  {1'b1,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b0,	1'b0,	ST_WAIT_MB};
        {ST_WAIT_MB,	1'b0,	1'bx,	1'b1}:tmp1265807652120  <=  {1'b1,	1'b0,	1'b1,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b0,	1'b0,	ST_REQ_M0};
        {ST_WAIT_MB,	1'b1,	1'b0,	1'b1}:tmp1265807652120  <=  {1'b1,	1'b0,	1'b1,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b0,	1'b0,	ST_REQ_M1};

        {ST_REQ_M0,	1'bx,	1'bx,	1'bx}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b0,	1'b1,	1'b0,	1'b0,	ST_WAIT_M0};

        {ST_WAIT_M0,	1'bx,	1'bx,	1'b0}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b0,	1'b1,	1'b0,	1'b0,	ST_WAIT_M0};
        {ST_WAIT_M0,	1'bx,	1'bx,	1'b1}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b0,	1'b0,	ST_REQ_MB};

        {ST_REQ_M1,	1'bx,	1'bx,	1'bx}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b0,	1'b0,	1'b0,	ST_WAIT_M1};

        {ST_WAIT_M1,	1'bx,	1'bx,	1'b0}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b0,	1'b0,	1'b0,	ST_WAIT_M1};
        {ST_WAIT_M1,	1'bx,	1'bx,	1'b1}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b1,	1'b0,	1'b0,	ST_REQ_MB};

        {ST_BOOTEND1,	1'bx,	1'bx,	1'bx}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b0,	1'b1,	ST_BOOTEND2};
        {ST_BOOTEND2,	1'bx,	1'bx,	1'bx}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b0,	1'b1,	ST_BOOTEND3};
        {ST_BOOTEND3,	1'bx,	1'bx,	1'bx}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b0,	1'b1,	ST_BOOTEND4};
        {ST_BOOTEND4,	1'bx,	1'bx,	1'bx}:tmp1265807652120  <=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b1,	1'b1,	ST_BOOTEND4};
       				default:tmp1265807652120  	<=  {1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b0,	1'b1,	1'b1,	1'b1,	1'b1,	1'b1,	ST_BOOTEND4};
    endcase
// This module was generated by xls2v on Wed Feb 10 22:14:12 GMT+09:00 2010.
endmodule

